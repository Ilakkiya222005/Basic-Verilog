module fourbit_twocom(